R0102 20296 20295 1
C0100 20296 20040 1
V0200 20295 20039 DC 10
= 19783 20039
- 20040 20039
.TRAN 20555 20554 TRAN 10 1
